`ifndef INCLUDE_SV
`define INCLUDE_SV
`include "transaction/item.sv"
`include "transaction/interface.sv"
`include "component/generator.sv"
`include "component/driver.sv"
`include "component/monitor.sv"
`include "component/scoreboard.sv"
`endif