package gcd_pkg;
  import uvm_pkg::*;
  `include "transaction/item.sv"
  `include "component/sequencer.sv"
  `include "component/generator.sv"
  `include "component/driver.sv"
  `include "component/monitor.sv"
  `include "component/scoreboard.sv"
  `include "component/agent.sv"
  `include "component/env.sv"
  `include "component/test.sv"
endpackage
